module MEM_WB_Latch ();

endmodule