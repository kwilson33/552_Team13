module ID_EX_Latch();

endmodule