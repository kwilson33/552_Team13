module Hazard_Detector ();


endmodule
