module EX_MEM_Latch ();

	input
	output

endmodule