module EX_MEM_Latch ();

endmodule